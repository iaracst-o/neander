module ula(
    input logic[7:0] ac,
    input logic [7:0] rdm,
    input logic [2:0] c,
    input logic [7:0] resul,
    output logic n,z
);


    
endmodule